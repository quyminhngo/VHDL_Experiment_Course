library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity BCDCounterSystem is
  port (
    resetn: in std_logic;
    pause: in std_logic
  );
end entity;

architecture RTL_BCDCounterSystem of BCDCounterSystem is
begin
    
    
end architecture;
